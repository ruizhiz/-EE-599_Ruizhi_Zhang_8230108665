module add(input [7:0] a, input [7:0] b, input [7:0] out);
	assign out = a + b;
endmodule
